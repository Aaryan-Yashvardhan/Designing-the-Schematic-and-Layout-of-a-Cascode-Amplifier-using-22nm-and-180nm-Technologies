magic
tech scmos
timestamp 1699270999
<< nwell >>
rect -97 114 117 115
rect -118 26 117 114
rect -118 -80 116 26
<< ntransistor >>
rect -87 -99 -55 -96
rect -25 -101 -23 -91
rect 21 -101 23 -91
rect 61 -101 63 -91
rect -25 -125 -23 -115
rect 21 -125 23 -115
rect 61 -125 63 -115
<< ptransistor >>
rect 37 10 42 19
rect -78 -23 -76 1
rect -37 -23 -35 1
rect -8 -13 4 -7
rect 37 -43 42 -34
<< ndiffusion >>
rect -95 -98 -94 -96
rect -90 -98 -87 -96
rect -95 -99 -87 -98
rect -55 -99 -51 -96
rect -35 -97 -25 -91
rect -35 -101 -33 -97
rect -29 -101 -25 -97
rect -23 -95 -18 -91
rect -14 -95 -12 -91
rect -23 -101 -12 -95
rect 10 -95 11 -91
rect 15 -95 21 -91
rect 10 -101 21 -95
rect 23 -97 33 -91
rect 23 -101 25 -97
rect 29 -101 33 -97
rect 51 -97 61 -91
rect 51 -101 54 -97
rect 58 -101 61 -97
rect 63 -93 66 -91
rect 70 -93 74 -91
rect 63 -101 74 -93
rect -34 -119 -33 -115
rect -29 -119 -25 -115
rect -34 -125 -25 -119
rect -23 -121 -11 -115
rect -23 -125 -16 -121
rect 10 -119 15 -115
rect 19 -119 21 -115
rect 10 -125 21 -119
rect 23 -121 33 -115
rect 23 -125 28 -121
rect 50 -121 61 -115
rect 50 -125 52 -121
rect 57 -125 61 -121
rect 63 -119 68 -115
rect 72 -119 73 -115
rect 63 -125 73 -119
<< pdiffusion >>
rect 31 14 37 19
rect 35 10 37 14
rect 42 15 44 19
rect 42 10 48 15
rect -97 -19 -78 1
rect -97 -23 -94 -19
rect -90 -23 -78 -19
rect -76 -1 -64 1
rect -76 -5 -68 -1
rect -76 -23 -64 -5
rect -49 -5 -48 1
rect -42 -5 -37 1
rect -49 -23 -37 -5
rect -35 -19 -23 1
rect -15 -11 -14 -7
rect -10 -11 -8 -7
rect -15 -13 -8 -11
rect 4 -9 11 -7
rect 4 -13 7 -9
rect -35 -23 -26 -19
rect 35 -38 37 -34
rect 31 -43 37 -38
rect 42 -37 48 -34
rect 42 -43 44 -37
<< ndcontact >>
rect -94 -98 -90 -94
rect -51 -100 -47 -96
rect -33 -101 -29 -97
rect -18 -95 -14 -91
rect 11 -95 15 -91
rect 25 -101 29 -97
rect 54 -101 58 -97
rect 66 -93 70 -89
rect -33 -119 -29 -115
rect -16 -125 -11 -121
rect 15 -119 19 -115
rect 28 -125 33 -121
rect 52 -125 57 -121
rect 68 -119 72 -115
<< pdcontact >>
rect 31 10 35 14
rect 44 15 48 19
rect -94 -23 -90 -19
rect -68 -5 -64 -1
rect -48 -5 -42 1
rect -14 -11 -10 -7
rect 7 -13 11 -9
rect -26 -23 -22 -19
rect 31 -38 35 -34
rect 44 -43 48 -37
<< psubstratepcontact >>
rect -48 -141 -41 -136
rect -27 -141 -20 -136
rect -8 -141 -1 -136
rect 14 -141 21 -136
rect 38 -141 45 -136
rect 61 -141 68 -136
<< nsubstratencontact >>
rect -89 43 -82 48
rect -54 44 -47 49
rect -21 44 -14 49
rect 4 44 11 49
rect 28 44 35 49
rect 49 44 56 49
<< polysilicon >>
rect 41 27 42 31
rect 37 19 42 27
rect -78 1 -76 2
rect -37 1 -35 6
rect -8 -7 4 6
rect 37 3 42 10
rect 37 -2 38 3
rect -8 -23 4 -13
rect -78 -25 -76 -23
rect -37 -25 -35 -23
rect -8 -27 0 -23
rect 37 -24 42 -22
rect 37 -29 38 -24
rect 37 -34 42 -29
rect 37 -48 42 -43
rect 37 -55 42 -52
rect -87 -90 -59 -86
rect -87 -96 -55 -90
rect -25 -91 -23 -90
rect 25 -87 59 -85
rect 21 -91 23 -89
rect 61 -91 63 -89
rect -87 -108 -55 -99
rect -25 -103 -23 -101
rect -25 -105 -7 -103
rect -3 -105 1 -103
rect 21 -102 23 -101
rect 5 -104 23 -102
rect 61 -104 63 -101
rect 21 -111 32 -109
rect 52 -109 53 -107
rect 52 -111 63 -109
rect -25 -113 -7 -111
rect -25 -115 -23 -113
rect -3 -113 2 -111
rect 6 -113 23 -111
rect 21 -115 23 -113
rect 61 -115 63 -111
rect -25 -129 -23 -125
rect 21 -129 23 -125
rect 61 -129 63 -125
<< polycontact >>
rect 37 27 41 31
rect -78 2 -74 6
rect 38 -2 42 3
rect -78 -29 -74 -25
rect -39 -29 -35 -25
rect 0 -27 4 -23
rect 38 -29 42 -24
rect 37 -52 42 -48
rect -59 -90 -55 -86
rect -27 -90 -23 -86
rect 21 -89 25 -85
rect 59 -89 63 -85
rect -7 -105 -3 -101
rect 1 -105 5 -101
rect 32 -111 36 -107
rect 47 -111 52 -107
rect -7 -115 -3 -111
rect 2 -115 6 -111
<< metal1 >>
rect -93 49 62 50
rect -93 48 -54 49
rect -93 43 -89 48
rect -82 44 -54 48
rect -47 44 -21 49
rect -14 44 4 49
rect 11 44 28 49
rect 35 44 49 49
rect 56 44 62 49
rect -82 43 62 44
rect -93 42 62 43
rect -74 2 -68 6
rect -64 -5 -58 42
rect -48 1 -42 42
rect -14 -7 -10 42
rect 28 27 37 31
rect 44 19 48 42
rect -94 -80 -90 -23
rect -22 -23 -21 -19
rect -74 -29 -39 -25
rect -26 -80 -21 -23
rect 0 -47 4 -27
rect 7 -47 12 -13
rect 31 -34 35 10
rect 42 -2 68 3
rect 42 -29 53 -24
rect 63 -37 68 -2
rect 48 -43 69 -37
rect 0 -48 12 -47
rect 0 -51 37 -48
rect 7 -52 37 -51
rect -94 -83 -50 -80
rect -26 -83 -14 -80
rect -94 -94 -90 -83
rect -53 -86 -50 -83
rect -18 -84 -14 -83
rect 7 -82 12 -52
rect -55 -90 -27 -86
rect -18 -88 -4 -84
rect 7 -86 16 -82
rect -18 -91 -14 -88
rect -51 -135 -47 -100
rect -33 -115 -29 -101
rect -7 -101 -3 -88
rect 11 -91 15 -86
rect 25 -89 59 -85
rect 66 -89 70 -43
rect 1 -101 5 -94
rect 25 -105 28 -101
rect -7 -111 -3 -105
rect 15 -108 28 -105
rect 55 -105 59 -101
rect -7 -116 -3 -115
rect 2 -122 6 -115
rect 15 -115 19 -108
rect 36 -111 47 -107
rect 55 -108 71 -105
rect 68 -115 71 -108
rect -16 -135 -11 -125
rect 28 -135 33 -125
rect 52 -135 57 -125
rect -51 -136 77 -135
rect -51 -141 -48 -136
rect -41 -141 -27 -136
rect -20 -141 -8 -136
rect -1 -141 14 -136
rect 21 -141 38 -136
rect 45 -141 61 -136
rect 68 -141 77 -136
<< labels >>
rlabel metal1 -72 44 -65 46 1 VDD
rlabel metal1 4 -140 8 -137 1 GND
rlabel metal1 -72 3 -68 6 1 Vbiasp
rlabel metal1 2 -122 6 -119 1 Vbias4
rlabel metal1 1 -100 5 -97 1 Vbias3
rlabel metal1 49 -28 53 -25 1 Vbias2
rlabel metal1 30 28 34 31 1 Vbias1
<< end >>
